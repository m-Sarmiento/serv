localparam [3:0]
  CSR_MSCRATCH  = 4'b0000,
  CSR_MTVEC     = 4'b0001,
  CSR_MEPC      = 4'b0010,
  CSR_MTVAL     = 4'b0011,
  CSR_DCSR      = 4'b0100,
  CSR_DPC       = 4'b0101,
  CSR_DSCRATCH0 = 4'b0110,
  CSR_DSCRATCH1 = 4'b0111,
  CSR_MHARTID   = 4'b1000,
  CSR_MISA      = 4'b1001;
